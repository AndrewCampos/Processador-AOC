module memoria(dado, endereco, write, wclk, rclk, saida);

	input [31:0] dado;
	input [9:0] endereco;
	input write, wclk, rclk;
	output reg [31:0] saida;
	reg [31:0]ram[127:0];
	
	initial begin	
		
		// GCD
		ram[10'd0] = 32'b00000100000111110000000111001101;  // addi
		ram[10'd1] = 32'b01010100000000000000000000011011;  // jmp
		ram[10'd2] = 32'b01000011111101000000000000000001;  // str
		ram[10'd3] = 32'b01000011111101010000000000000010;  // str
		ram[10'd4] = 32'b01000111111000010000000000000010;  // ldr
		ram[10'd5] = 32'b00000100000000100000000000000000;  // addi
		ram[10'd6] = 32'b00101100010000010000000000001011;  // bne
		ram[10'd7] = 32'b01000111111001000000000000000001;  // ldr
		ram[10'd8] = 32'b00000100100111100000000000000000;  // addi
		ram[10'd9] = 32'b01011100000000000000000000000000;  // jst
		ram[10'd10] = 32'b01010100000000000000000000011010;   // jmp
		ram[10'd11] = 32'b01000111111001010000000000000010;   // ldr
		ram[10'd12] = 32'b00000100101101000000000000000000;   // addi
		ram[10'd13] = 32'b01000111111001100000000000000001;   // ldr
		ram[10'd14] = 32'b01000111111001110000000000000001;   // ldr
		ram[10'd15] = 32'b01000111111010000000000000000010;   // ldr
		ram[10'd16] = 32'b00000000111010000100100000000011;   // div
		ram[10'd17] = 32'b01000111111010100000000000000010;   // ldr
		ram[10'd18] = 32'b00000001001010100101100000000010;   // mult
		ram[10'd19] = 32'b00000000110010110110000000000001;   // sub
		ram[10'd20] = 32'b00000101100101010000000000000000;   // addi
		ram[10'd21] = 32'b00000111111111110000000000000010;   // addi
		ram[10'd22] = 32'b01011000000000000000000000000010;   // jal
		ram[10'd23] = 32'b00001011111111110000000000000010;   // subi
		ram[10'd24] = 32'b00000111110111100000000000000000;   // addi
		ram[10'd25] = 32'b01011100000000000000000000000000;   // jst
		ram[10'd26] = 32'b01011100000000000000000000000000;   // jst
		ram[10'd27] = 32'b01000111111011010000000000000001;   // ldr
		ram[10'd28] = 32'b01001100000111100000000000000000;   // in
		ram[10'd29] = 32'b00000111110011010000000000000000;   // addi
		ram[10'd30] = 32'b01000011111011010000000000000001;   // str
		ram[10'd31] = 32'b01000111111011100000000000000010;   // ldr
		ram[10'd32] = 32'b01001100000111100000000000000000;   // in
		ram[10'd33] = 32'b00000111110011100000000000000000;   // addi
		ram[10'd34] = 32'b01000011111011100000000000000010;   // str
		ram[10'd35] = 32'b00000111110101000000000000000000;   // addi
		ram[10'd36] = 32'b01010100000000000000000000100101;   // jmp
		ram[10'd37] = 32'b01001000000000000000000000000000;   // hlt
		
			
			
	end 
	always @ (posedge wclk)
	begin
		if (write == 1'b1)
			ram[endereco] <= dado;
	end
	
always @ (negedge rclk) saida <= ram[endereco];
	
endmodule
